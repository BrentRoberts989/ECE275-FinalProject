/*
*
*/
module paddle(paddleMove, )
	